/*
 * CODER: Luis Fernando Rodriguez Gtz
 * DATE: 14/Ago/2023
 * PROJECT: 
 */

`ifndef DIGITALTUBE_MUX_PKG_SV
    `define DIGITALTUBE_MUX_PKG_SV
package digitalTube_mux_pkg;
    /** Parameters*/
    /*  */
    localparam clkFreq_FPGA = 27_000_000;
    
    localparam clkFreq_TargetHz = 10_000;
 
endpackage: digitalTube_mux_pkg
`endif