/*
 * CODER: Luis Fernando Rodriguez Gtz
 * DATE: 14/Ago/2023
 * PROJECT: 
 */
 
 import common_pkg::*;
 
 module digitalTube
(
    /** INPUT*/
    input data2display_t display_data,
    /** OUTPUT*/
    output digital_tube_t digital_tube_enable
);
	
/* Obtain the numbers necesary to ignite each display */ 
always_comb 
begin

end 
endmodule
